`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 12/07/2024 11:14:38 PM
// Design Name: 
// Module Name: Diff_sub_mod
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module Diff_sub_mod();

    //subtractor subtractor1(result window1 frame1)
    //subtractor subtractor2(result window1 frame1) ect
    
    
    //add abs functions or code that into the subtractors idk



endmodule
