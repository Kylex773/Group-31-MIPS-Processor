`timescale 1ns / 1ps

////////////////////////////////////////////////////////////////////////////////
// ECE369A - Computer Architecture
// Laboratory 1
// Module - ProgramCounter_tb.v
// Description - Test the 'ProgramCounter.v' module.
////////////////////////////////////////////////////////////////////////////////

module ProgramCounter_tb(); 

	reg [31:0] Address;
	reg Reset, Clk;

	wire [31:0] PCResult;

    ProgramCounter u0(
        .Address(Address), 
        .PCResult(PCResult), 
        .Reset(Reset), 
        .Clk(Clk)
    );

	initial begin
		Clk <= 1'b0;
		forever #15 Clk <= ~Clk;
	end

	initial begin
	
    /* Please fill in the implementation here... */
    Reset <=1;
    #80;
    
    Reset <=0;
    
    Address<=20;
	#30;
	
	Address<=2;
	#30;

	Address<=50;
	#30;
	
	Address<=100;
	#30;
    end
	


endmodule

