`timescale 1ns / 1ps

////////////////////////////////////////////////////////////////////////////////
// ECE369A - Computer Architecture
// Laboratory  
// Module - PCAdder.v
// Description - 32-Bit program counter (PC) adder.
// 
// INPUTS:-
// PCResult: 32-Bit input port.
// 
// OUTPUTS:-
// PCAddResult: 32-Bit output port.
//
// FUNCTIONALITY:-
// Design an incrementor (or a hard-wired ADD ALU whose first input is from the 
// PC, and whose second input is a hard-wired 4) that computes the current 
// PC + 4. The result should always be an increment of the signal 'PCResult' by 
// 4 (i.e., PCAddResult = PCResult + 4).
////////////////////////////////////////////////////////////////////////////////

module PCAdder(PCResult, PCAddResult);

    input [31:0] PCResult;

    output reg [31:0] PCAddResult;

    /* Please fill in the implementation here... */
    
    always @(PCResult, PCAddResult) begin
        PCAddResult <= PCResult + 4;
        
    end
endmodule
    
    
    /*`timescale 1ns / 1ps

//A + B + Cin gives S and Co where Co is Carry-out
module Adder_12bits(A, B, Cin, S, Co);
    
    input [11:0] A, B;
    input Cin;
    output reg [11:0] S;
    output reg Co;
    
    //write your code here
    always @(A,B,Cin) begin
    
        {Co, S} <= A + B + Cin;
    
    end

endmodule
*/



